module present_tb ();

`ifdef PERIOD
  parameter time period = `PERIOD ;
`else
  parameter time period = 40ns ;
`endif


import present_pkg::*;

logic clk = 0;
logic nrst = 0;
logic start = 0;
wire eoc;
logic [63:0] plaintext = '0;
logic [127:0]key = '0;
wire  [63:0] ciphertext;

logic [63:0] D[0:4] = '{{64{1'b0}},{64{1'b0}},{64{1'b1}},{64{1'b1}}, 64'h0123456789abcdef};
logic [127:0]K[0:4] = '{{128{1'b0}},{128{1'b1}},{128{1'b0}},{128{1'b1}}, 128'h0123456789abcdef0123456789abcdef};

`ifdef USE_VAMS_WRAPPER
bit energy_measurement ;
real measured_energy ;

breadboard dut    (
		     .clk(clk),
                    .nrst(nrst),
                    .start(start),
                    .eoc(eoc),
                    .plaintext(plaintext),
                    .key(key),
                    .ciphertext(ciphertext),
                    .energy_measurement(energy_measurement),
                    .measured_energy(measured_energy)
		   );
`else
present_v0 dut    (
                    .clk(clk),
                    .nrst(nrst),
                    .start(start),
                    .eoc(eoc),
                    .plaintext(plaintext),
                    .key(key),
                    .ciphertext(ciphertext)
               );
`endif
// clock
always #(period/2) clk = !clk;

// Files for vcd and info
`ifndef vcdfilename
`define  vcdfilename  "../results/present_v0.vcd"
`endif
`ifndef vcdinfofile
`define  vcdinfofile  "../results/present_v0_vcd_info.tcl"
`endif
// File for results and measurements
`define  resultfile "../results/results.dat"
integer fr ; // pointer to the file containing infos for VCD
integer fres ; // pointer to the file containing simulation results

initial
   $display("---- clock period %p", period);

initial
begin
    $display("Unrolled %3d times", ROUNDS_PER_CYCLE);
end

initial
begin
   int i;
   fres = $fopen(`resultfile,"w") ;
   $timeformat(-12,0,"",6) ;
   $fdisplay(fres, "Testing the 128bit   version of present");
   $fdisplay(fres, "Unrolled %3d times", ROUNDS_PER_CYCLE);
   $fdisplay(fres,"---- clock period %tps", period);

   `ifdef DUMP_VCD
     $dumpfile(`vcdfilename) ;
     $dumpvars(0,present_tb.dut) ;
   //  $dumpoff;
     fr = $fopen(`vcdinfofile,"w") ;
     $fwrite(fr,"# Generated by \"sim\" process\n# Time in ps\n");
     $timeformat(-12,0,"",20) ;
     $fwrite(fr,"set vcd_start %0t\n",$realtime);
   `endif
   plaintext = $random();
   key = $random();

   // reset
   repeat(4) @(posedge clk);
   #(period/2) ;
   nrst = 1;
   `ifdef USE_VAMS_WRAPPER
    energy_measurement = 1'b1 ;
   `endif
   repeat(4) @(posedge clk);
   // start of test
   for (i=0; i<5; i++)
   begin
      @(posedge  clk);
      #(period/2) ;
      plaintext = D[i];
      key       = K[i];
      start = 1;
      @(posedge clk);
      #(period/2) ;
      start = 0;
      forever @(posedge clk)
      begin
         if (eoc) break;
      end
      assert (ciphertext == PCrypt(D[i],K[i]))
      begin
         $info ("%x (+) %x -> %x",D[i], K[i], ciphertext);
	 $fdisplay(fres,"%x (+) %x -> %x",D[i], K[i], ciphertext) ;
      end
      else
      begin
         $fatal (0, "%x (+) %x -> %x !!error!! should be %x",D[i], K[i], ciphertext,PCrypt(D[i],K[i]));
      end
   end
   $fdisplay(fres,"----- End of simulation -----");
   @(posedge  clk);

   `ifdef USE_VAMS_WRAPPER
    energy_measurement = 1'b0 ;
   `endif
   `ifdef DUMP_VCD
     $timeformat(-12,0,"",20) ;
     $fwrite(fr,"set vcd_stop %0t\n",$realtime);
     $fclose(fr);
   `endif
    @(posedge  clk);
   `ifdef USE_VAMS_WRAPPER
      $fdisplay(fres,"Measured energy: %fpJ",measured_energy*1.0e12) ;
   `endif
   $fclose(fr) ;
   $fclose(fres);
   $finish();
end

endmodule
